**.subckt vco_2-4GHz_tb
V1 vctl 0 vctl
Vdd net1 0 vdd
xvco net1 Ip In Qp Qn NCp NCn FBp FBn vctl 0 vco_2-4GHz
**** begin user architecture code


.param temp=125.000000
.temp 125.000000

.save v(ip) v(in) v(vctl) i(vdd)

.include sky130_fd_pr/cells/rf_pfet_01v8_lvt/sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35.spice
.lib sky130_fd_pr/models/sky130.lib.spice lh
.tran 0.01n 10n uic
.param vdd=1.800000
.param vctl=1.800000


**** end user architecture code
**.ends

* expanding   symbol:  vco_2-4GHz/vco_2-4GHz.sym # of pins=11

.subckt vco_2-4GHz  VDD ph1_p ph1_n ph2_p ph2_n ph3_p ph3_n ph4_p ph4_n CTL GND
*.ipin CTL
*.iopin VDD
*.iopin GND
*.opin ph3_p
*.opin ph3_n
*.opin ph4_p
*.opin ph4_n
*.opin ph2_p
*.opin ph2_n
*.opin ph1_p
*.opin ph1_n
x1 VDD net2 net1 net7 net8 GND CTL vco_2-4Ghz_delaycell
x2 VDD net4 net3 net2 net1 GND CTL vco_2-4Ghz_delaycell
x3 VDD net6 net5 net4 net3 GND CTL vco_2-4Ghz_delaycell
x4 VDD net8 net7 net6 net5 GND CTL vco_2-4Ghz_delaycell
x5 VDD ph1_p ph1_n net1 net2 GND rf_bufferdiff
x6 VDD ph2_p ph2_n net3 net4 GND rf_bufferdiff
x7 VDD ph3_p ph3_n net5 net6 GND rf_bufferdiff
x8 VDD ph4_p ph4_n net7 net8 GND rf_bufferdiff
I0 GND GND pulse(1000n 0 0 400p 100p 100p 10 20 0)
.ends


* expanding   symbol:  vco_2-4GHz_delaycell/vco_2-4Ghz_delaycell.sym # of pins=7

.subckt vco_2-4Ghz_delaycell  VDD OUTn OUTp Pn Pp GND CTL
*.ipin Pp
*.ipin Pn
*.opin OUTn
*.opin OUTp
*.iopin VDD
*.iopin GND
*.ipin CTL
XXMprimpos OUTp Pp GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 m=3
XXMcrossneg OUTn OUTp GND GND sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 m=1
XXMctlneg OUTn CTL VDD VDD sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 m=1
XXMctlpos OUTp CTL VDD VDD sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 m=1
XXMcrosspos OUTp OUTn GND GND sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 m=1
XXMprimneg OUTn Pn GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 m=3
XXMctlpos1 net2 GND VDD VDD sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 m=1
XXMctlneg1 net1 GND VDD VDD sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 m=1
XXMctlpos2 OUTp GND net2 VDD sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 m=1
XXMctlneg2 OUTn GND net1 VDD sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 m=1
.ends


* expanding   symbol:  rf_bufferdiff/rf_bufferdiff.sym # of pins=6

.subckt rf_bufferdiff  vdd out_n out_p in_p in_n vss
*.iopin vdd
*.iopin vss
*.ipin in_p
*.ipin in_n
*.opin out_n
*.opin out_p
XXMdiffp out_n in_p vss vss sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 m=1
XXMdiffn out_p in_n vss vss sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 m=1
XRn vdd out_n vss sky130_fd_pr__res_xhigh_po_2p85 m=1
XRp vdd out_p vss sky130_fd_pr__res_xhigh_po_2p85 m=1
.ends

.end
