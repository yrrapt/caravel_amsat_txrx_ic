module user_project_wrapper(
            inout     vssd1,
            inout     vccd1,
            inout     vssd2,
            inout     vccd2,
            in        la_data_in[0],
            in        la_data_in[1],
            in        la_data_in[2],
            in        la_data_in[3],
            in        la_data_in[4],
            in        la_data_in[5],
            in        la_data_in[6],
            in        la_data_in[7],
            in        la_data_in[8],
            in        la_data_in[9],
            in        la_data_in[10],
            in        la_data_in[11],
            in        la_data_in[12],
            in        la_data_in[13],
            in        la_data_in[14],
            in        la_data_in[15],
            in        la_data_in[16],
            in        la_data_in[17],
            in        la_data_in[18],
            in        la_data_in[19],
            in        la_data_in[20],
            in        la_data_in[21],
            in        la_data_in[22],
            in        la_data_in[23],
            in        la_data_in[24],
            in        la_data_in[25],
            in        la_data_in[26],
            in        la_data_in[27],
            in        la_data_in[28],
            in        la_data_in[29],
            in        la_data_in[95],
            in        la_data_in[94],
            in        la_data_in[93],
            in        la_data_in[92],
            in        la_data_in[91],
            in        la_data_in[90],
            in        la_data_in[89],
            in        la_data_in[88],
            in        la_data_in[87],
            in        la_data_in[86],
            in        la_data_in[85],
            in        la_data_in[84],
            in        la_data_in[83],
            in        la_data_in[82],
            in        la_data_in[81],
            in        la_data_in[80],
            in        la_data_in[79],
            in        la_data_in[78],
            inout     analog_io[0],
            inout     analog_io[1],
            inout     analog_io[2],
            inout     analog_io[3],
            inout     analog_io[4],
            inout     analog_io[5],
            inout     analog_io[6],
            inout     analog_io[7],
            inout     analog_io[8],
            inout     analog_io[9],
            inout     analog_io[10],
            inout     analog_io[11],
            inout     analog_io[12],
            inout     analog_io[13],
            inout     analog_io[14],
            inout     analog_io[15],
            inout     analog_io[16],
            inout     analog_io[17],
            inout     analog_io[18],
            inout     analog_io[19],
            inout     analog_io[20],
            inout     analog_io[21],
            inout     analog_io[24],
            inout     analog_io[25],
            inout     analog_io[26],
            inout     analog_io[27],
            inout     analog_io[28],
            inout     analog_io[29],
            inout     analog_io[30]
    );


      fake fake ();



endmodule
